//Define a uvm environment class named apb_env
`ifndef apb_environment
`define apb_environment
`include "uvm_macros.svh"
import uvm_pkg::*;
import apb_pkg::*;

class apb_env extends uvm_env;
  
  //register the class with uvm factory
	`uvm_component_utils(apb_env)

	//	Component Members
	apb_master_agent  master_agent;
	apb_scoreboard    apb_scb;
	apb_env_config 	  apb_env_cfg;
  //virtual interface for apb interface
	virtual apb_if  vif;
  
  //constructor for the class
  function new(string name = "apb_env", uvm_component parent = null);
    //call the base class constructor
	  super.new(name, parent);
  endfunction
  
  //Build phase - construct agents, virtual sequencer and get virtual interface handle
  function void build_phase(uvm_phase phase);
	  super.build_phase(phase);
    //create an instance of the master agnet
  	master_agent = apb_master_agent::type_id::create("master_agent", this);
	if(apb_env_cfg ==null) begin
		uvm_config_db#(apb_env_config)::get(null,"","apb_env_config",apb_env_cfg);
	end
	if(apb_env_cfg.has_scoreboard) begin
		apb_scb =apb_scoreboard::type_id::create("apb_scb",this);
	end
    //create an instance of the slave agent
  	if (!uvm_config_db#(virtual apb_if)::get(null, "", "apb_vif", vif)) begin
		  `uvm_fatal(get_full_name(), "No virtual interface specified for env")
	  end		
  endfunction
  
  //connect phase
  function void connect_phase(uvm_phase phase);
    super.connect_phase(phase);
   // uvm_config_db#(apb_master_sequencer)::set(this,"*","master_seqr",master_agent.m_sequencer);
    //uvm_config_db#(apb_slave_sequencer)::set(this,"*","slave_seqr",slave_agent.m_sequencer);	
	if(apb_env_cfg.has_scoreboard) begin
  		master_agent.m_apb_master_monitor.ap.connect(apb_scb.ap_mntr2scb);
		master_agent.m_apb_master_driver.drv2scb.connect(apb_scb.ap_drv2scb);
	end
  endfunction
  
  //print topology
  function void end_of_elaboration_phase(uvm_phase phase);
    uvm_top.print_topology();
  endfunction
  
endclass  //end of the class
`endif
